`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/11/28 15:30:45
// Design Name: 
// Module Name: DMUX_32
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module decoder_32(
    input [4:0] waddr,
    input we,
    output reg [31:0] ena_d
    );
    always @(*)
           begin
              if(we == 0)
                ena_d=32'b0000_0000_0000_0000_0000_0000_0000_0000;
              else
              begin
               case(waddr)
                 5'd0: ena_d =  32'b0000_0000_0000_0000_0000_0000_0000_0001;
                 5'd1: ena_d =  32'b0000_0000_0000_0000_0000_0000_0000_0010;
                 5'd2: ena_d =  32'b0000_0000_0000_0000_0000_0000_0000_0100;
                 5'd3: ena_d =  32'b0000_0000_0000_0000_0000_0000_0000_1000;
                 5'd4: ena_d =  32'b0000_0000_0000_0000_0000_0000_0001_0000;
                 5'd5: ena_d =  32'b0000_0000_0000_0000_0000_0000_0010_0000;
                 5'd6: ena_d =  32'b0000_0000_0000_0000_0000_0000_0100_0000;
                 5'd7: ena_d =  32'b0000_0000_0000_0000_0000_0000_1000_0000;
                 5'd8: ena_d =  32'b0000_0000_0000_0000_0000_0001_0000_0000;
                 5'd9: ena_d =  32'b0000_0000_0000_0000_0000_0010_0000_0000;
                 5'd10: ena_d = 32'b0000_0000_0000_0000_0000_0100_0000_0000;
                 5'd11: ena_d = 32'b0000_0000_0000_0000_0000_1000_0000_0000;
                 5'd12: ena_d = 32'b0000_0000_0000_0000_0001_0000_0000_0000;
                 5'd13: ena_d = 32'b0000_0000_0000_0000_0010_0000_0000_0000;
                 5'd14: ena_d = 32'b0000_0000_0000_0000_0100_0000_0000_0000;
                 5'd15: ena_d = 32'b0000_0000_0000_0000_1000_0000_0000_0000;
                 5'd16: ena_d = 32'b0000_0000_0000_0001_0000_0000_0000_0000;
                 5'd17: ena_d = 32'b0000_0000_0000_0010_0000_0000_0000_0000;
                 5'd18: ena_d = 32'b0000_0000_0000_0100_0000_0000_0000_0000;
                 5'd19: ena_d = 32'b0000_0000_0000_1000_0000_0000_0000_0000;
                 5'd20: ena_d = 32'b0000_0000_0001_0000_0000_0000_0000_0000;
                 5'd21: ena_d = 32'b0000_0000_0010_0000_0000_0000_0000_0000;
                 5'd22: ena_d = 32'b0000_0000_0100_0000_0000_0000_0000_0000;
                 5'd23: ena_d = 32'b0000_0000_1000_0000_0000_0000_0000_0000;
                 5'd24: ena_d = 32'b0000_0001_0000_0000_0000_0000_0000_0000;
                 5'd25: ena_d = 32'b0000_0010_0000_0000_0000_0000_0000_0000;
                 5'd26: ena_d = 32'b0000_0100_0000_0000_0000_0000_0000_0000;
                 5'd27: ena_d = 32'b0000_1000_0000_0000_0000_0000_0000_0000;
                 5'd28: ena_d = 32'b0001_0000_0000_0000_0000_0000_0000_0000;
                 5'd29: ena_d = 32'b0010_0000_0000_0000_0000_0000_0000_0000;
                 5'd30: ena_d = 32'b0100_0000_0000_0000_0000_0000_0000_0000;
                 5'd31: ena_d = 32'b1000_0000_0000_0000_0000_0000_0000_0000;
                 
               endcase
               end
            end
endmodule
